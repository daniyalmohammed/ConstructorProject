0
0 0 0 0 0 r h 0 B 17 B
0 0 0 0 0 r h 4 B 15 B
0 0 0 0 0 r h 2 B 20 B
0 0 0 0 0 r h 6 B 10 B
3 11 2 9 0 9 1 12 4 8 1 3 4 6 0 10 0 8 1 11 1 4 3 4 4 3 5 7 2 5 0 10 2 2 3 5 2 6
4
