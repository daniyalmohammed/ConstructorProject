1
10 9 13 9 13 r 0 2 4 8 16 24 h 0 B 4 T 10 B 22 H
1 1 1 1 0 r 70 h 15 H 53 B
0 0 0 0 0 r 36 41 h 27 B 34 T
2 3 3 4 6 r 43 45 47 54 55 60 h 30 H 37 B 42 H
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
7
